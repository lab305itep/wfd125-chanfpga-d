localparam VERSION = 32'h00000201;